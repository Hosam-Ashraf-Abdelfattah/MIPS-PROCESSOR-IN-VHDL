library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_arith.ALL;
--use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all; 


--library UNISIM;
--use UNISIM.VComponents.all;

entity fetchingg is
			port(
			clk:in std_logic ;
			reset:in std_logic ;
			pc_src_control:in std_logic:='0' ;
			pc_pranch_src :in std_logic_vector (31 downto 0);
								
  				
  			RD_ADDR		: out	STD_LOGIC_VECTOR (4 downto 0);
			RS_ADDR		: out	STD_LOGIC_VECTOR (4 downto 0);
			RT_ADDR		: out	STD_LOGIC_VECTOR (4 downto 0);
			ofset			: out	STD_LOGIC_VECTOR (15 downto 0);
			funct		: out	STD_LOGIC_VECTOR (5 downto 0);
			READ_ADDR2 :out std_logic_vector (31 downto 0);
			re_fitch	: in	STD_LOGIC:='0';
			INST_simulation : out std_logic_vector (31 downto 0);
			opcode		: out	STD_LOGIC_VECTOR (5 downto 0));
			
		
end fetchingg;

architecture Behavioral of fetchingg is


 signal READ_ADDR	: 	STD_LOGIC_VECTOR (31 downto 0);
 signal INST		: 	STD_LOGIC_VECTOR (31 downto 0);
begin


	
	
	process (clk,reset)
	begin
	if reset='1' then
	READ_ADDR <="00000000000000000000000000000000";
	
--	elsif(rising_edge(clk))then
--		if re_fitch='0' then
--			if pc_src_control = '0' then
--				READ_ADDR <= READ_ADDR + 4;
--			else 
--				READ_ADDR <= pc_pranch_src;
--			end if;
--		else
--						READ_ADDR <= READ_ADDR;
--		end if;
--	end if;
	elsif(rising_edge(clk))then
		if re_fitch='0' and pc_src_control = '0' then
			
				READ_ADDR <= READ_ADDR + 4;
		elsif re_fitch='0' and pc_src_control = '1' then
				READ_ADDR <= pc_pranch_src;
			
		else
						READ_ADDR <= READ_ADDR;
		end if;
	end if;
	end process;
	READ_ADDR2 <= READ_ADDR + 4;
----------------------------------------------------------------------------	
	process (READ_ADDR)
	begin

		case READ_ADDR is
			when "00000000000000000000000000000000" => 
				INST <= "01010001010000100010001000100000";
			when "00000000000000000000000000000100" => 
				INST <= "10001100010100001000000000100010";
			when "00000000000000000000000000001000" => 
				INST <= "00110000110000100000000000100010";
			when "00000000000000000000000000001100" => 
				INST <= "00101110001101010000000000100010";
			when "00000000000000000000000000010000" => 
				INST <= "00010101110001100001011000100010";
			when "00000000000000000000000000010100" => 
				INST <= "00010100100100010001100100100000";
			when "00000000000000000000000000011000" => 
				INST <= "00101000101001000010000000100010";
			when "00000000000000000000000000011100" => 
				INST <= "00010000100000100000100000100010";
			when "00000000000000000000000000100000" => 
				INST <= "00110000100001000000100100100010";
			when "00000000000000000000000000100100" => 
				INST <= "00100000010000000000000000100010";
			when "00000000000000000000000000101000" => 
				INST <= "10010000011000110010000000100000";
			when "00000000000000000000000000101100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000000110000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000000110100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000000111000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000000111100" => 
				INST <= "00000000100010110010000000100010";
			when "00000000000000000000000001000000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000001000100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000001001000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000001001100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000001010000" => 
				INST <= "00000000100000000100000000101010";
			when "00000000000000000000000001010100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000001011000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000001011100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000001100000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000001100100" => 
				INST <= "00010001000000010000000000001000";
			when "00000000000000000000000001101000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000001101100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000001110000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000001110100" => 
				INST <= "00000001100001010110000000100101";
			when "00000000000000000000000001111000" => 
				INST <= "00010000000000000000000000000100";
			when "00000000000000000000000001111100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000010000000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000010000100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000010001000" => 
				INST <= "00000000011000110010000000100000";
			when "00000000000000000000000010001100" => 
				INST <= "00000000110000010011000000100000";
			when "00000000000000000000000010010000" => 
				INST <= "00000000101001010010100000100000";
			when "00000000000000000000000010010100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000010011000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000010011100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000010100000" => 
				INST <= "00000000110001110100000000101010";
			when "00000000000000000000000010100100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000010101000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000010101100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000010110000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000010110100" => 
				INST <= "00010001000000011111111111010111";
			when others => 
				INST <= "11111111111111111111111111111111";
				
		end case;
----------------------------------------------------------------
	end process;
	process(INST)
	begin
	funct<=INST(5 downto 0);
	RD_ADDR<=INST(15 downto 11);
	RT_ADDR<=INST(20 downto 16);
	RS_ADDR<=INST(25 downto 21);
	opcode<=INST(31 downto 26);
	ofset<=INST(15 downto 0);
	INST_simulation<=READ_ADDR;
	end process;
	
	


end Behavioral;